/* minimig_defines.v */
/* 2012, rok.krajnc@gmail.com */

`define MINIMIG_ALTERA
