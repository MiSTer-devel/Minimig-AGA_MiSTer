// minimig version constants

localparam [7:0] BETA_FLAG = 8'd1;  // BETA / RELEASE flag
localparam [7:0] MAJOR_VER = 8'd1;  // major version number
localparam [7:0] MINOR_VER = 8'd2;  // minor version number
localparam [7:0] SEPARATOR = 8'd0;  // separator (should be set to 0)

